module I2C_AV_Config(
	// Host Side
	o_I2C_END,
	iCLK,
	iRST_N,
	iVOL,

	// I2C Side
	I2C_SCLK,
	I2C_SDAT
);

	// Host Side
	input iCLK;
	input iRST_N;
	input [6:0] iVOL;

	// I2C Side
	output I2C_SCLK;
	inout I2C_SDAT;
	output o_I2C_END ;

	// Internal Registers/Wires
	reg	[15:0] mI2C_CLK_DIV;
	reg	[23:0] mI2C_DATA;
	reg mI2C_CTRL_CLK;
	reg	mI2C_GO;
	wire mI2C_END;
	wire mI2C_ACK;
	reg	[15:0] LUT_DATA;
	reg	[3:0] LUT_INDEX;
	reg	[1:0] mSetup_ST;
	reg o_I2C_END;

	// Clock Setting
	parameter CLK_Freq = 50000000; // 50 MHz
	parameter I2C_Freq = 20000; // 20 KHz

	// LUT Data Number
	parameter LUT_SIZE = 12;

	//	Audio Data Index
	parameter Dummy_DATA = 0;
	parameter REG_REST = 1;
	parameter SET_LIN_L	= 2;
	parameter SET_LIN_R	= 3;
	parameter SET_HEAD_L = 4;
	parameter SET_HEAD_R = 5;
	parameter A_PATH_CTRL =	6;
	parameter D_PATH_CTRL =	7;
	parameter POWER_ON = 8;
	parameter SET_FORMAT = 9;
	parameter SAMPLE_CTRL =	10;
	parameter SET_ACTIVE = 11;

	// I2C Control Clock
	always @(posedge iCLK or negedge iRST_N) begin
		if (!iRST_N) begin
			mI2C_CTRL_CLK <= 0;
			mI2C_CLK_DIV <= 0;
		end else begin
			if (mI2C_CLK_DIV < (CLK_Freq/I2C_Freq))
				mI2C_CLK_DIV <=	mI2C_CLK_DIV+1;
			else begin
				mI2C_CLK_DIV <=	0;
				mI2C_CTRL_CLK <= ~mI2C_CTRL_CLK;
			end
		end
	end

	I2C_Controller u0(
		.CLOCK(mI2C_CTRL_CLK), // Controller Work Clock
		.I2C_SCLK(I2C_SCLK), //	I2C CLOCK
		.I2C_SDAT(I2C_SDAT), //	I2C DATA
		.I2C_DATA(mI2C_DATA), // DATA:[SLAVE_ADDR,SUB_ADDR,DATA]
		.GO(mI2C_GO),  // GO transfor
		.END(mI2C_END), // END transfor 
		.ACK(mI2C_ACK), // ACK
		.RESET(iRST_N)
	);

	// Config Control
	always @(posedge mI2C_CTRL_CLK or negedge iRST_N) begin
		if (!iRST_N) begin
			LUT_INDEX <= 0;
			mSetup_ST <= 0;
			mI2C_GO <= 0;
		end else begin
			if (LUT_INDEX < LUT_SIZE) begin
				o_I2C_END <= 0 ;

				case(mSetup_ST)
					0: begin
						mI2C_DATA <= {8'h34,LUT_DATA};
						mI2C_GO <= 1;
						mSetup_ST <= 1;
					end
					1: begin
						if (mI2C_END) begin
							if (!mI2C_ACK)
								mSetup_ST <= 2;
							else
								mSetup_ST <= 0;							
								mI2C_GO <= 0;
						end
					end
					2: begin
						LUT_INDEX <= LUT_INDEX + 1;
						mSetup_ST <= 0;
					end
				endcase
			end else begin
				o_I2C_END <= 1;
			end
		end
	end

	// Config Data LUT
	always begin
		case(LUT_INDEX) // Audio Config Data
			Dummy_DATA: LUT_DATA <= 16'h0000;
			REG_REST: LUT_DATA <= 16'h1E00;
			SET_LIN_L: LUT_DATA <= 16'h001A;
			SET_LIN_R: LUT_DATA	<= 16'h021A;
			SET_HEAD_L: LUT_DATA <=	{8'h04, 1'b1, iVOL};
			SET_HEAD_R: LUT_DATA <=	{8'h06, 1'b1, iVOL};
			A_PATH_CTRL: LUT_DATA <= 16'h08F8;
			D_PATH_CTRL: LUT_DATA <= 16'h0A06;
			POWER_ON: LUT_DATA <= 16'h0C00;
			SET_FORMAT: LUT_DATA <=	16'h0E01;
			SAMPLE_CTRL: LUT_DATA <= 16'h1002;
			SET_ACTIVE:	LUT_DATA <=	16'h1201;
			default: LUT_DATA <= 16'h0000;
		endcase
	end

endmodule
