module wave_gen_sin(
	input [7:0] ramp,
	input clk,
	output [15:0] music_o
);

	reg [15:0] music;
	always @(ramp[7:0]) begin
		case(ramp[7:0])
			 0: music = 16'h0000;
			 1: music = 16'h0349;
			 2: music = 16'h038D;
			 3: music = 16'h008D;
			 4: music = 16'hFD0B;
			 5: music = 16'hFC41;
			 6: music = 16'hFEE9;
			 7: music = 16'h0291;
			 8: music = 16'h03DD;
			 9: music = 16'h019C;
			10: music = 16'hFDE0;
			11: music = 16'hFC18;
			12: music = 16'hFDE7;
			13: music = 16'h01A4;
			14: music = 16'h03DF;
			15: music = 16'h028A;
			16: music = 16'hFEE0;
			17: music = 16'hFC3F;
			18: music = 16'hFD11;
			19: music = 16'h0096;
			20: music = 16'h0391;
			21: music = 16'h0345;
			22: music = 16'hFFF7;
			23: music = 16'hFCB2;
			24: music = 16'hFC76;
			25: music = 16'hFF7C;
			26: music = 16'h02FB;
			27: music = 16'h03BC;
			28: music = 16'h010F;
			29: music = 16'hFD68;
			30: music = 16'hFC24;
			31: music = 16'hFE6C;
			32: music = 16'h0227;
			33: music = 16'h03E8;
			34: music = 16'h0211;
			35: music = 16'hFE54;
			36: music = 16'hFC20;
			37: music = 16'hFD7C;
			38: music = 16'h0128;
			39: music = 16'h03C4;
			40: music = 16'h02E9;
			41: music = 16'hFF61;
			42: music = 16'hFC6B;
			43: music = 16'hFCC0;
			44: music = 16'h0012;
			45: music = 16'h0353;
			46: music = 16'h0386;
			47: music = 16'h007C;
			48: music = 16'hFD00;
			49: music = 16'hFC46;
			50: music = 16'hFEFA;
			51: music = 16'h029E;
			52: music = 16'h03DB;
			53: music = 16'h018C;
			54: music = 16'hFDD1;
			55: music = 16'hFC18;
			56: music = 16'hFDF6;
			57: music = 16'h01B4;
			58: music = 16'h03E1;
			59: music = 16'h027D;
			60: music = 16'hFECF;
			61: music = 16'hFC3A;
			62: music = 16'hFD1D;
			63: music = 16'h00A7;
			64: music = 16'h0398;
			65: music = 16'h033B;
			66: music = 16'hFFE5;
			67: music = 16'hFCA8;
			68: music = 16'hFC7E;
			69: music = 16'hFF8D;
			70: music = 16'h0306;
			71: music = 16'h03B7;
			72: music = 16'h00FE;
			73: music = 16'hFD5B;
			74: music = 16'hFC27;
			75: music = 16'hFE7C;
			76: music = 16'h0236;
			77: music = 16'h03E8;
			78: music = 16'h0202;
			79: music = 16'hFE44;
			80: music = 16'hFC1E;
			81: music = 16'hFD8A;
			82: music = 16'h0139;
			83: music = 16'h03C8;
			84: music = 16'h02DD;
			85: music = 16'hFF50;
			86: music = 16'hFC65;
			87: music = 16'hFCCA;
			88: music = 16'h0023;
			89: music = 16'h035C;
			90: music = 16'h037E;
			91: music = 16'h006A;
			92: music = 16'hFCF5;
			93: music = 16'hFC4C;
			94: music = 16'hFF0B;
			95: music = 16'h02AB;
			96: music = 16'h03D8;
			97: music = 16'h017C;
			98: music = 16'hFDC3;
			99: music = 16'hFC19;
		   100: music = 16'hFE06;
		   101: music = 16'h01C4;
		   102: music = 16'h03E3;
		   103: music = 16'h026F;
		   104: music = 16'hFEBE;
		   105: music = 16'hFC35;
		   106: music = 16'hFD29;
		   107: music = 16'h00B9;
		   108: music = 16'h039F;
		   109: music = 16'h0331;
		   110: music = 16'hFFD4;
		   111: music = 16'hFC9F;
		   112: music = 16'hFC86;
		   113: music = 16'hFF9F;
		   114: music = 16'h0311;
		   115: music = 16'h03B1;
		   116: music = 16'h00ED;
		   117: music = 16'hFD4E;
		   118: music = 16'hFC2A;
		   119: music = 16'hFE8D;
		   120: music = 16'h0245;
		   121: music = 16'h03E7;
		   122: music = 16'h01F3;
		   123: music = 16'hFE34;
		   124: music = 16'hFC1C;
		   125: music = 16'hFD98;
		   126: music = 16'h014A;
		   127: music = 16'h03CD;
		   128: music = 16'h02D1;
		   129: music = 16'hFF3F;
		   130: music = 16'hFC5E;
		   131: music = 16'hFCD4;
		   132: music = 16'h0035;
		   133: music = 16'h0365;
		   134: music = 16'h0376;
		   135: music = 16'h0058;
		   136: music = 16'hFCEA;
		   137: music = 16'hFC51;
		   138: music = 16'hFF1C;
		   139: music = 16'h02B8;
		   140: music = 16'h03D4;
		   141: music = 16'h016B;
		   142: music = 16'hFDB4;
		   143: music = 16'hFC1A;
		   144: music = 16'hFE15;
		   145: music = 16'h01D4;
		   146: music = 16'h03E4;
		   147: music = 16'h0261;
		   148: music = 16'hFEAE;
		   149: music = 16'hFC31;
		   150: music = 16'hFD35;
		   151: music = 16'h00CA;
		   152: music = 16'h03A5;
		   153: music = 16'h0326;
		   154: music = 16'hFFC2;
		   155: music = 16'hFC97;
		   156: music = 16'hFC8E;
		   157: music = 16'hFFB0;
		endcase
	end
	
	assign music_o = music;

endmodule
