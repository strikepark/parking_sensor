module hex_7seg(
	input [3:0] cs,
	input [3:0] ds,
	input [3:0] s,
	input [3:0] das,

	output reg [6:0] seg0,
	output reg [6:0] seg1,
	output reg [6:0] seg2,
	output reg [6:0] seg3
);

	always @(cs[3:0]) begin
		case (cs[3:0])
			4'b0000: seg0 <= 7'b1_00_00_00;
			4'b0001: seg0 <= 7'b1_11_10_01;
			4'b0010: seg0 <= 7'b0_10_01_00;
			4'b0011: seg0 <= 7'b0_11_00_00;
			4'b0100: seg0 <= 7'b0_01_10_01;
			4'b0101: seg0 <= 7'b0_01_00_10;
			4'b0110: seg0 <= 7'b0_00_00_10;
			4'b0111: seg0 <= 7'b1_11_10_00;
			4'b1000: seg0 <= 7'b0_00_00_00;
			4'b1001: seg0 <= 7'b0_01_00_00;
			default: seg0 <= 7'b1_11_11_11;
		endcase
	end

	always @(ds[3:0]) begin
		case (ds[3:0])
			4'b0000: seg1 <= 7'b1_00_00_00;
			4'b0001: seg1 <= 7'b1_11_10_01;
			4'b0010: seg1 <= 7'b0_10_01_00;
			4'b0011: seg1 <= 7'b0_11_00_00;
			4'b0100: seg1 <= 7'b0_01_10_01;
			4'b0101: seg1 <= 7'b0_01_00_10;
			4'b0110: seg1 <= 7'b0_00_00_10;
			4'b0111: seg1 <= 7'b1_11_10_00;
			4'b1000: seg1 <= 7'b0_00_00_00;
			4'b1001: seg1 <= 7'b0_01_00_00;
			default: seg1 <= 7'b1_11_11_11;
		endcase
	end

	always @(s[3:0]) begin
		case (s[3:0])
			4'b0000: seg2 <= 7'b1_00_00_00;
			4'b0001: seg2 <= 7'b1_11_10_01;
			4'b0010: seg2 <= 7'b0_10_01_00;
			4'b0011: seg2 <= 7'b0_11_00_00;
			4'b0100: seg2 <= 7'b0_01_10_01;
			4'b0101: seg2 <= 7'b0_01_00_10;
			4'b0110: seg2 <= 7'b0_00_00_10;
			4'b0111: seg2 <= 7'b1_11_10_00;
			4'b1000: seg2 <= 7'b0_00_00_00;
			4'b1001: seg2 <= 7'b0_01_00_00;
			default: seg2 <= 7'b1_11_11_11;
		endcase
	end

	always @(das[3:0]) begin
		case (das[3:0])
			4'b0000: seg3 <= 7'b1_00_00_00;
			4'b0001: seg3 <= 7'b1_11_10_01;
			4'b0010: seg3 <= 7'b0_10_01_00;
			4'b0011: seg3 <= 7'b0_11_00_00;
			4'b0100: seg3 <= 7'b0_01_10_01;
			4'b0101: seg3 <= 7'b0_01_00_10;
			4'b0110: seg3 <= 7'b0_00_00_10;
			4'b0111: seg3 <= 7'b1_11_10_00;
			4'b1000: seg3 <= 7'b0_00_00_00;
			4'b1001: seg3 <= 7'b0_01_00_00;
			default: seg3 <= 7'b1_11_11_11;
		endcase
	end

endmodule
